** sch_path: /home/swati/work/xschem/OP2.sch
**.subckt OP2
R1 vn1 vn2 5k m=1
R2 vn2 vout 5k m=1
C1 vin vn1 4.7u m=1
V1 vin GND AC 1 sin(0 1m 1e3 0 0 0)
V2 net1 GND 1.5
x2 vout net1 vn2 GND opamp_model
**** begin user architecture code



* ngspice commands
.control
OP
save all
write Complete_ckt.raw
set appendwrite
Ac DEC 100 1 10e6
plot vdb(vout)
plot v(vout)
plot phase(vout)
MEAS AC gain_db MAX vdb(vout) FROM=1 TO=10e6
LET vm3db = gain_db-3.0
print vm3db
MEAS AC fzero WHEN vdb(vout)=vm3db RISE=1
MEAS AC fpole WHEN vdb(vout)=vm3db FALL=1
** phase measurement
LET phase_deg = cph(vout)*180/PI
MEAS AC phase_zero FIND phase_deg AT=fzero
MEAS AC phase_pole FIND phase_deg AT=fpole
MEAS AC phase_mid FIND phase_deg AT=fmid
** MEAS fero fpole using phase
LET phase_zero_ph = phase_mid - 45
MEAS AC fzero_ph WHEN phase_deg=phase_zero_ph
.endc
.end


**** end user architecture code
**.ends

* expanding   symbol:  opamp_model.sym # of pins=4
** sym_path: /home/swati/work/xschem/opamp_model.sym
** sch_path: /home/swati/work/xschem/opamp_model.sch
.subckt opamp_model vop vip vim vom
*.iopin vop
*.iopin vom
*.iopin vip
*.iopin vim
E1 vop vom vip vim 1000
.ends

.GLOBAL GND
.end
