** sch_path: /home/swati/work/xschem/op.sch
**.subckt op
V3 vnmic GND 0 AC 1
R4 vnmic vn1 380 m=1
C4 vn1 vn2 4.7u m=1
R5 vn2 net1 4.7k m=1
R6 net1 vout 300k m=1
C5 net1 vout 27p m=1
C6 vout GND 1p m=1
V4 net2 GND 1.5
**** begin user architecture code



* ngspice commands
.control
op
save all
write mictest.raw
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
