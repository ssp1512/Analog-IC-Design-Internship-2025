** sch_path: /home/swati/work/xschem/mictestop.sch
**.subckt mictestop
V1 vnmic GND 0 AC 1
R1 vnmic vn1 380 m=1
C1 vn1 vn2 4.7u m=1
R2 vn2 net2 4.7k m=1
R3 net2 net3 300k m=1
C2 net2 net3 27p m=1
C3 net3 GND 1p m=1
V2 net1 GND 1.5
x1 net3 net2 net1 GND opamp_model
**** begin user architecture code



* ngspice commands
.control
OP
save all
write Complete_ckt.raw
set appendwrite
Ac DEC 100 1 10e6
plot vdb(vout)
plot v(vout)
plot phase(vout)
MEAS AC gain_db MAX vdb(vout) FROM=1 TO=10e6
LET vm3db = gain_db-3.0
print vm3db
MEAS AC fzero WHEN vdb(vout)=vm3db RISE=1
MEAS AC fpole WHEN vdb(vout)=vm3db FALL=1
** phase measurement
LET phase_deg = cph(vout)*180/PI
MEAS AC phase_zero FIND phase_deg AT=fzero
MEAS AC phase_pole FIND phase_deg AT=fpole
MEAS AC phase_mid FIND phase_deg AT=fmid
** MEAS fero fpole using phase
LET phase_zero_ph = phase_mid - 45
MEAS AC fzero_ph WHEN phase_deg=phase_zero_ph
.endc
.end


**** end user architecture code
**.ends

* expanding   symbol:  opamp_model.sym # of pins=4
** sym_path: /home/swati/work/xschem/opamp_model.sym
** sch_path: /home/swati/work/xschem/opamp_model.sch
.subckt opamp_model vop vip vim vom
*.iopin vop
*.iopin vom
*.iopin vip
*.iopin vim
E1 vop vom vip vim 1000
.ends

.GLOBAL GND
.end
