** sch_path: /home/swati/work/xschem/oplowsch
**.subckt oplowsch
E1 net1 net4 vn2 net3 1000
E2 vout GND net2 net4 1
R1 net1 net2 1k m=1
C1 net2 net4 160n m=1
R2 vn1 vn2 5k m=1
R3 vn2 vout 5k m=1
C2 vin vn1 4.7u m=1
V1 vin GND 0 AC 1
V2 net3 GND 1.5
**** begin user architecture code



* ngspice commands
.control
.OP
AC DEC 100 1 10e6
plot v(vout)
.ENDC


**** end user architecture code
**.ends
.GLOBAL GND
.end
