** sch_path: /home/swati/work/xschem/op4.sch
**.subckt op4
R1 vn1 vn2 5k m=1
R2 vn2 vout 5k m=1
C1 vin vn1 4.7u m=1
V1 vin GND AC 1 sin(0 1m 1e3 0 0 0)
V2 net1 GND 1.5
x1 vout net1 vn2 GND op3
**** begin user architecture code



* ngspice commands
.control
OP
save all
write Complete_ckt.raw
set appendwrite
Ac DEC 100 1 10e6
plot vdb(vout)
plot v(vout)
plot phase(vout)
MEAS AC gain_db MAX vdb(vout) FROM=1 TO=10e6
LET vm3db = gain_db-3.0
print vm3db
MEAS AC fzero WHEN vdb(vout)=vm3db RISE=1
MEAS AC fpole WHEN vdb(vout)=vm3db FALL=1
** phase measurement
LET phase_deg = cph(vout)*180/PI
MEAS AC phase_zero FIND phase_deg AT=fzero
MEAS AC phase_pole FIND phase_deg AT=fpole
MEAS AC phase_mid FIND phase_deg AT=fmid
** MEAS fero fpole using phase
LET phase_zero_ph = phase_mid - 45
MEAS AC fzero_ph WHEN phase_deg=phase_zero_ph
.endc
.end


**** end user architecture code
**.ends

* expanding   symbol:  op3.sym # of pins=4
** sym_path: /home/swati/work/xschem/op3.sym
** sch_path: /home/swati/work/xschem/op3.sch
.subckt op3 vop vinp vinm vom
*.iopin vinp
*.iopin vinm
*.iopin vop
*.iopin vom
E1 net1 net3 vinp vinm 3
E2 vop vom net2 net3 3
R1 net1 net2 1k m=1
C1 net2 net3 160n m=1
.ends

.GLOBAL GND
.end
