** sch_path: /home/swati/work/xschem/lowapss.sch
**.subckt lowapss vop vom
*.iopin vop
*.iopin vom
R1 vn1 vn2 5k m=1
R2 vn2 vout 5k m=1
C1 vin vn1 4.7u m=1
V1 vin GND 0 AC 1
V2 net4 GND 1.5
E1 net1 net3 vn2 net4 1000
E2 vop vom net2 net3 1000
R3 net1 net2 1k m=1
C2 net2 net3 160n m=1
**** begin user architecture code



* ngspice commands
.control
.op
AC DEC 100 1 10e6
plot v(vout)
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
